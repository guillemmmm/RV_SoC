/********1*********2*********3*********4*********5*********6*********7*********8
* File : spi_defines.vh
*_______________________________________________________________________________
*
* Revision history
*
* Name          Date        Observations
* ------------------------------------------------------------------------------
* -            01/02/2022   First version.
* ------------------------------------------------------------------------------
*_______________________________________________________________________________
*
* Description
* SPI master macro definition file
*_______________________________________________________________________________

* (c) Copyright Universitat de Barcelona, 2022
*
*********1*********2*********3*********4*********5*********6*********7*********/
// SPI MASTER REGISTERS ADDRESS
`define SPI_CTRL   2'h0
`define SPI_BUFFER 2'h1
`define SPI_CONFIG 2'h2
`define SPI_SSELEC 2'h3
